library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rect_renderer is
  port (
    clk : in std_logic;
    reset : in boolean;
    go : in boolean;
  );
end entity;

architecture rtl of rect_renderer is

begin



end architecture;
